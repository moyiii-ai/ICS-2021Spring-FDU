`include "common.svh"