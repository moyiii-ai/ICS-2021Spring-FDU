`include "common.svh"

module decode (

);

endmodule