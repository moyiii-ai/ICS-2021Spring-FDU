`ifndef __ICODE_SVH__
`define __ICODE_SVH__

`define LUI 6'b001111