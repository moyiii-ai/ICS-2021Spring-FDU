`include "common.svh"

module hazard(

);

endmodule